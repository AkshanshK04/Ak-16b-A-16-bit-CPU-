module cpu_tb;
    reg clk;
    reg rst;

    // Instantiate CPU
    cpu_top dut(
        .clk(clk),
        .rst(rst)
    );

    // Clock generation - 10ns period (100MHz)
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    // Test sequence
    initial begin
        // Dump waveforms
        $dumpfile("cpu.vcd");
        $dumpvars(0, cpu_tb);

        // Display register values
        $display("\n=== AK-16 CPU Simulation Started ===\n");
        $monitor("T=%0t | PC=%h Instr=%h Op=%h | R1=%h R2=%h R3=%h R4=%h | MemW=%b RegW=%b", 
                 $time, dut.pc, dut.instr, dut.opcode,
                 dut.u_rf.regs[1], dut.u_rf.regs[2], 
                 dut.u_rf.regs[3], dut.u_rf.regs[4],
                 dut.mem_write, dut.reg_write);
        // Reset sequence
        rst = 1;
        #15;
        rst = 0;
        
        // Run for sufficient time
        #500;
        
        // Display final register state
        $display("\n=== Final Register State ===");
        $display("R0=%h R1=%h R2=%h R3=%h", 
                 dut.u_rf.regs[0], dut.u_rf.regs[1],
                 dut.u_rf.regs[2], dut.u_rf.regs[3]);
        $display("R4=%h R5=%h R6=%h R7=%h",
                 dut.u_rf.regs[4], dut.u_rf.regs[5],
                 dut.u_rf.regs[6], dut.u_rf.regs[7]);
        $display("R8=%h R9=%h RA=%h RB=%h",
                 dut.u_rf.regs[8], dut.u_rf.regs[9],
                 dut.u_rf.regs[10], dut.u_rf.regs[11]);
        $display("RC=%h RD=%h RE=%h RF=%h",
                 dut.u_rf.regs[12], dut.u_rf.regs[13],
                 dut.u_rf.regs[14], dut.u_rf.regs[15]);
        
        //to view memory contents
        $display("\n=== Memory Contents ===");
        $display("mem[0]=%h mem[1]=%h mem[2]=%h mem[3]=%h",
                 dut.u_dmem.mem[0], dut.u_dmem.mem[1],
                 dut.u_dmem.mem[2], dut.u_dmem.mem[3]);

        $finish;
    end
    //Watchdog for HALT detection
    always @(posedge clk) begin
        if (dut.instr == 16'hF00 && !rst ) begin
            #20;
            $display("\n=== HALT Instruction Detected at PC=%h===", dut.pc);
            $display("\n=== All Registers (Hex/Dec) ===");
            $display("R0 = %04h (%5d)    R1 = %04h (%5d)", 
                     dut.u_rf.regs[0], dut.u_rf.regs[0],
                     dut.u_rf.regs[1], dut.u_rf.regs[1]);
            $display("R2 = %04h (%5d)    R3 = %04h (%5d)", 
                     dut.u_rf.regs[2], dut.u_rf.regs[2],
                     dut.u_rf.regs[3], dut.u_rf.regs[3]);
            $display("R4 = %04h (%5d)    R5 = %04h (%5d)", 
                     dut.u_rf.regs[4], dut.u_rf.regs[4],
                     dut.u_rf.regs[5], $signed(dut.u_rf.regs[5]));
            $display("R6 = %04h (%5d)    R7 = %04h (%5d)", 
                     dut.u_rf.regs[6], dut.u_rf.regs[6],
                     dut.u_rf.regs[7], dut.u_rf.regs[7]);
            $display("R8 = %04h (%5d)    R9 = %04h (%5d)", 
                     dut.u_rf.regs[8], dut.u_rf.regs[8],
                     dut.u_rf.regs[9], dut.u_rf.regs[9]);
            $display("RA = %04h (%5d)    RB = %04h (%5d)", 
                     dut.u_rf.regs[10], dut.u_rf.regs[10],
                     dut.u_rf.regs[11], dut.u_rf.regs[11]);
            $display("RC = %04h (%5d)    RD = %04h (%5d)", 
                     dut.u_rf.regs[12], dut.u_rf.regs[12],
                     dut.u_rf.regs[13], dut.u_rf.regs[13]);
            $display("RE = %04h (%5d)    RF = %04h (%5d)", 
                     dut.u_rf.regs[14], dut.u_rf.regs[14],
                     dut.u_rf.regs[15], dut.u_rf.regs[15]);
            #10;
            $finish;
        end
    end
endmodule